**.subckt reram_example
.inc sky130_fd_pr_reram__reram_cell.spice

V1 TE 0 PWL (0 0 0.25u 1.4 0.5u 0 0.75u -1.4 1.0u 0.0)
XR0 TE 0 sky130_fd_pr_reram__reram_cell Tfilament_0=3.3e-9

.tran 0.1n 1.5u

.end